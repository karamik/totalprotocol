// TOTAL Protocol Sentinel Core v.8.0 Hardware Interface
